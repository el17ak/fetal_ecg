package fsm_fastica;


endpackage
