module invert_mat #(
	parameter SIZE_A = 8,
	parameter SIZE_B = 8,
	parameter N_BITS = 22
)
(
	input reading matrix [SIZE_A][SIZE_B],
	output reading out[SIZE_A][SIZE_B]
);

endmodule
