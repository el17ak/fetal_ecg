module eigenvalue_decomposition #(
	parameter SIZE_N = 8
	
)
(
	input integer mat[SIZE_N][SIZE_N],
	output integer eigenvector_mat[SIZE_N][SIZE_N],
	output integer eigenvalues[SIZE_N]
);



endmodule
