module uart_tx #(
	parameter SIZE_A,
	parameter SIZE_B,
	parameter N_BITS
)
(
	input clk,
	input logic[N_BITS-1:0] matrix[SIZE_A][SIZE_B]
);

	

endmodule
