package fsm_eigenloop;

	typedef enum{
		INITIALISATION_EIGEN,
		WAIT_EIGEN,
		RECURSION_EIGEN,
		CONVERGENCE_EIGEN,
		FINISHED_EIGEN,
		XXX_EIGEN
	} state_eigenloop;

endpackage
