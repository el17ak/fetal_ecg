module bluetooth_tx(

);

endmodule
