module invert_mat #(
	parameter SIZE_A = 8,
	parameter SIZE_B = 8
)
(
	input integer matrix [SIZE_A][SIZE_B],
	output integer out[SIZE_A][SIZE_B]
);

endmodule
