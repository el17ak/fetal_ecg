module whiten(
	input logic clk,
	input logic[7:0][7:0] matrix
);

//D * D'

endmodule
