module uart_rx(
	input clk
);


endmodule
