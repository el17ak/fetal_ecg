module trigger_while(

)
(
	input logic trigger,
	input 
);